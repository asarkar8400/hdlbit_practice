module top_module ( input a, input b, output out );
    mod_a instance2 ( a, b, out );
endmodule
